----------------------------------------------------------------------------------
-- Company:  Gruppe 2 - Semesterprojekt 2014

-- Module Name:    		main - Behavioral
-- Module description:  

-- Change date		Engineer 
-- 06-03-2014 		ALB
--
--
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

----------------------------------------------------------------------------------

entity main is
end main;

architecture Behavioral of main is

begin


end Behavioral;

